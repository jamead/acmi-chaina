------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version : 3.6
--  \   \         Application : 7 Series FPGAs Transceivers Wizard 
--  /   /         Filename : kria_comm_support.vhd
-- /___/   /\      
-- \   \  /  \ 
--  \___\/\___\
--
--  Description : This module instantiates the modules required for
--                reset and initialisation of the Transceiver
--
-- Module kria_comm_support
-- Generated by Xilinx 7 Series FPGAs Transceivers Wizard
-- 
-- 
-- (c) Copyright 2010-2012 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;
--***********************************Entity Declaration************************

entity kria_comm_support is
generic
(
    EXAMPLE_SIM_GTRESET_SPEEDUP             : string    := "TRUE";     -- simulation setting for GT SecureIP model
    STABLE_CLOCK_PERIOD                     : integer   := 10  

);
port
(
    SOFT_RESET_TX_IN                        : in   std_logic;
    SOFT_RESET_RX_IN                        : in   std_logic;
    DONT_RESET_ON_DATA_ERROR_IN             : in   std_logic;
    Q0_CLK0_GTREFCLK_PAD_N_IN               : in   std_logic;
    Q0_CLK0_GTREFCLK_PAD_P_IN               : in   std_logic;
    refclk_out                              : out  std_logic;

    GT0_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_DATA_VALID_IN                       : in   std_logic;
    GT0_TX_MMCM_LOCK_OUT                    : out  std_logic;
    GT0_RX_MMCM_LOCK_OUT                    : out  std_logic;
 
    GT0_TXUSRCLK_OUT                        : out  std_logic;
    GT0_TXUSRCLK2_OUT                       : out  std_logic;
    GT0_RXUSRCLK_OUT                        : out  std_logic;
    GT0_RXUSRCLK2_OUT                       : out  std_logic;

    --_________________________________________________________________________
    --GT0  (X0Y0)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt0_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt0_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt0_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt0_drpen_in                            : in   std_logic;
    gt0_drprdy_out                          : out  std_logic;
    gt0_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt0_eyescanreset_in                     : in   std_logic;
    gt0_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt0_eyescandataerror_out                : out  std_logic;
    gt0_eyescantrigger_in                   : in   std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt0_rxdata_out                          : out  std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt0_rxchariscomma_out                   : out  std_logic_vector(3 downto 0);
    gt0_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    gt0_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt0_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt0_gtprxn_in                           : in   std_logic;
    gt0_gtprxp_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt0_rxcommadet_out                      : out  std_logic;
    gt0_rxmcommaalignen_in                  : in   std_logic;
    gt0_rxpcommaalignen_in                  : in   std_logic;
    ------------ Receive Ports - RX Decision Feedback Equalizer(DFE) -----------
    gt0_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt0_rxlpmhfhold_in                      : in   std_logic;
    gt0_rxlpmlfhold_in                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt0_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt0_gtrxreset_in                        : in   std_logic;
    gt0_rxlpmreset_in                       : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt0_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt0_gttxreset_in                        : in   std_logic;
    gt0_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt0_txdata_in                           : in   std_logic_vector(31 downto 0);
    ------------------ Transmit Ports - TX 8B/10B Encoder Ports ----------------
    gt0_txcharisk_in                        : in   std_logic_vector(3 downto 0);
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    gt0_gtptxn_out                          : out  std_logic;
    gt0_gtptxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt0_txoutclkfabric_out                  : out  std_logic;
    gt0_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt0_txresetdone_out                     : out  std_logic;

    --____________________________COMMON PORTS________________________________
   GT0_PLL0RESET_OUT  : out std_logic;
         GT0_PLL0OUTCLK_OUT  : out std_logic;
         GT0_PLL0OUTREFCLK_OUT  : out std_logic;
         GT0_PLL0LOCK_OUT  : out std_logic;
         GT0_PLL0REFCLKLOST_OUT  : out std_logic;    
         GT0_PLL1OUTCLK_OUT  : out std_logic;
         GT0_PLL1OUTREFCLK_OUT  : out std_logic;
       sysclk_in        : in std_logic

);

end kria_comm_support;
    
architecture RTL of kria_comm_support is
attribute DowngradeIPIdentifiedWarnings: string;
attribute DowngradeIPIdentifiedWarnings of RTL : architecture is "yes";

--**************************Component Declarations*****************************

component kria_comm
 
port
(
    SYSCLK_IN                               : in   std_logic;
    SOFT_RESET_TX_IN                        : in   std_logic;
    SOFT_RESET_RX_IN                        : in   std_logic;
    DONT_RESET_ON_DATA_ERROR_IN             : in   std_logic;
    GT0_DRP_BUSY_OUT                        : out  std_logic;
    GT0_TX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_RX_FSM_RESET_DONE_OUT               : out  std_logic;
    GT0_DATA_VALID_IN                       : in   std_logic;
    GT0_TX_MMCM_LOCK_IN                     : in   std_logic;
    GT0_TX_MMCM_RESET_OUT                   : out  std_logic;
    GT0_RX_MMCM_LOCK_IN                     : in   std_logic;
    GT0_RX_MMCM_RESET_OUT                   : out  std_logic;

    --_________________________________________________________________________
    --GT0  (X0Y0)
    --____________________________CHANNEL PORTS________________________________
    ---------------------------- Channel - DRP Ports  --------------------------
    gt0_drpaddr_in                          : in   std_logic_vector(8 downto 0);
    gt0_drpclk_in                           : in   std_logic;
    gt0_drpdi_in                            : in   std_logic_vector(15 downto 0);
    gt0_drpdo_out                           : out  std_logic_vector(15 downto 0);
    gt0_drpen_in                            : in   std_logic;
    gt0_drprdy_out                          : out  std_logic;
    gt0_drpwe_in                            : in   std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    gt0_eyescanreset_in                     : in   std_logic;
    gt0_rxuserrdy_in                        : in   std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    gt0_eyescandataerror_out                : out  std_logic;
    gt0_eyescantrigger_in                   : in   std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    gt0_rxdata_out                          : out  std_logic_vector(31 downto 0);
    gt0_rxusrclk_in                         : in   std_logic;
    gt0_rxusrclk2_in                        : in   std_logic;
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    gt0_rxchariscomma_out                   : out  std_logic_vector(3 downto 0);
    gt0_rxcharisk_out                       : out  std_logic_vector(3 downto 0);
    gt0_rxdisperr_out                       : out  std_logic_vector(3 downto 0);
    gt0_rxnotintable_out                    : out  std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    gt0_gtprxn_in                           : in   std_logic;
    gt0_gtprxp_in                           : in   std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    gt0_rxcommadet_out                      : out  std_logic;
    gt0_rxmcommaalignen_in                  : in   std_logic;
    gt0_rxpcommaalignen_in                  : in   std_logic;
    ------------ Receive Ports - RX Decision Feedback Equalizer(DFE) -----------
    gt0_dmonitorout_out                     : out  std_logic_vector(14 downto 0);
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    gt0_rxlpmhfhold_in                      : in   std_logic;
    gt0_rxlpmlfhold_in                      : in   std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    gt0_rxoutclk_out                        : out  std_logic;
    gt0_rxoutclkfabric_out                  : out  std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    gt0_gtrxreset_in                        : in   std_logic;
    gt0_rxlpmreset_in                       : in   std_logic;
    ----------------- Receive Ports - RX Polarity Control Ports ----------------
    gt0_rxpolarity_in                       : in   std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    gt0_rxresetdone_out                     : out  std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    gt0_gttxreset_in                        : in   std_logic;
    gt0_txuserrdy_in                        : in   std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    gt0_txdata_in                           : in   std_logic_vector(31 downto 0);
    gt0_txusrclk_in                         : in   std_logic;
    gt0_txusrclk2_in                        : in   std_logic;
    ------------------ Transmit Ports - TX 8B/10B Encoder Ports ----------------
    gt0_txcharisk_in                        : in   std_logic_vector(3 downto 0);
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    gt0_gtptxn_out                          : out  std_logic;
    gt0_gtptxp_out                          : out  std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    gt0_txoutclk_out                        : out  std_logic;
    gt0_txoutclkfabric_out                  : out  std_logic;
    gt0_txoutclkpcs_out                     : out  std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    gt0_txresetdone_out                     : out  std_logic;


    --____________________________COMMON PORTS________________________________
         GT0_PLL0OUTCLK_IN  : in std_logic;
         GT0_PLL0OUTREFCLK_IN  : in std_logic;
   GT0_PLL0RESET_OUT  : out std_logic;
         GT0_PLL0LOCK_IN  : in std_logic;
         GT0_PLL0REFCLKLOST_IN  : in std_logic;    
         GT0_PLL1OUTCLK_IN  : in std_logic;
         GT0_PLL1OUTREFCLK_IN  : in std_logic

);

end component;

component kria_comm_common_reset  
generic
(
      STABLE_CLOCK_PERIOD      : integer := 8        -- Period of the stable clock driving this state-machine, unit is [ns]
   );
port
   (    
      STABLE_CLOCK             : in std_logic;             --Stable Clock, either a stable clock from the PCB
      SOFT_RESET               : in std_logic;               --User Reset, can be pulled any time
      COMMON_RESET             : out std_logic  --Reset QPLL
   );
end component;

component kria_comm_common 
generic
(
    -- Simulation attributes
    WRAPPER_SIM_GTRESET_SPEEDUP     : string     :=  "FALSE" ;       -- Set to "TRUE" to speed up sim reset
    SIM_PLL0REFCLK_SEL              :bit_vector  := "001";
    SIM_PLL1REFCLK_SEL              :bit_vector  := "001"
 
);
port
(
    PLL0OUTCLK_OUT       : out std_logic;
    PLL0OUTREFCLK_OUT    : out std_logic;
    PLL0LOCK_OUT         : out std_logic;
    PLL0LOCKDETCLK_IN    : in std_logic;
    PLL0REFCLKLOST_OUT   : out std_logic;    
    PLL0RESET_IN         : in std_logic;
    PLL0REFCLKSEL_IN     : in std_logic_vector(2 downto 0);
    PLL0PD_IN            : in std_logic;
    PLL1OUTCLK_OUT       : out std_logic;
    PLL1OUTREFCLK_OUT    : out std_logic;
    GTREFCLK1_IN         : in std_logic;
    GTREFCLK0_IN         : in std_logic

);

end component;

component kria_comm_cpll_railing
  Generic(
           USE_BUFG       : integer := 0
);
port 
(   
        cpll_reset_out : out std_logic;
         cpll_pd_out : out std_logic;
         refclk_out : out std_logic;
        
         refclk_in : in std_logic

);
end component;
component kria_comm_GT_USRCLK_SOURCE 
port
(
 
    GT0_TXUSRCLK_OUT             : out std_logic;
    GT0_TXUSRCLK2_OUT            : out std_logic;
    GT0_TXOUTCLK_IN              : in  std_logic;
    GT0_TXCLK_LOCK_OUT           : out std_logic;
    GT0_TX_MMCM_RESET_IN         : in std_logic;
    GT0_RXUSRCLK_OUT             : out std_logic;
    GT0_RXUSRCLK2_OUT            : out std_logic;
    GT0_RXOUTCLK_IN              : in  std_logic;
    GT0_RXCLK_LOCK_OUT           : out std_logic;
    GT0_RX_MMCM_RESET_IN         : in std_logic;
    Q0_CLK0_GTREFCLK_PAD_N_IN               : in   std_logic;
    Q0_CLK0_GTREFCLK_PAD_P_IN               : in   std_logic;
    Q0_CLK0_GTREFCLK_OUT                    : out  std_logic
);
end component;

--***********************************Parameter Declarations********************

    constant DLY : time := 1 ns;

--************************** Register Declarations ****************************

    signal   gt0_txfsmresetdone_i            : std_logic;
signal   gt0_rxfsmresetdone_i            : std_logic;
    signal   gt0_txfsmresetdone_r            : std_logic;
    signal   gt0_txfsmresetdone_r2           : std_logic;
signal   gt0_rxresetdone_r               : std_logic;
signal   gt0_rxresetdone_r2              : std_logic;
signal   gt0_rxresetdone_r3              : std_logic;


signal   reset_pulse                     : std_logic_vector(3 downto 0);
    signal   reset_counter  :   unsigned(5 downto 0) := "000000";

--**************************** Wire Declarations ******************************
    -------------------------- GT Wrapper Wires ------------------------------
    --________________________________________________________________________
    --________________________________________________________________________
    --GT0  (X0Y0)

    ---------------------------- Channel - DRP Ports  --------------------------
    signal  gt0_drpaddr_i                   : std_logic_vector(8 downto 0);
    signal  gt0_drpdi_i                     : std_logic_vector(15 downto 0);
    signal  gt0_drpdo_i                     : std_logic_vector(15 downto 0);
    signal  gt0_drpen_i                     : std_logic;
    signal  gt0_drprdy_i                    : std_logic;
    signal  gt0_drpwe_i                     : std_logic;
    ------------------------ GTPE2_CHANNEL Clocking Ports ----------------------
    signal  gt0_pll0clk_i                   : std_logic;
    signal  gt0_pll0refclk_i                : std_logic;
    signal  gt0_pll1clk_i                   : std_logic;
    signal  gt0_pll1refclk_i                : std_logic;
    --------------------- RX Initialization and Reset Ports --------------------
    signal  gt0_eyescanreset_i              : std_logic;
    signal  gt0_rxuserrdy_i                 : std_logic;
    -------------------------- RX Margin Analysis Ports ------------------------
    signal  gt0_eyescandataerror_i          : std_logic;
    signal  gt0_eyescantrigger_i            : std_logic;
    ------------------ Receive Ports - FPGA RX Interface Ports -----------------
    signal  gt0_rxdata_i                    : std_logic_vector(31 downto 0);
    ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
    signal  gt0_rxchariscomma_i             : std_logic_vector(3 downto 0);
    signal  gt0_rxcharisk_i                 : std_logic_vector(3 downto 0);
    signal  gt0_rxdisperr_i                 : std_logic_vector(3 downto 0);
    signal  gt0_rxnotintable_i              : std_logic_vector(3 downto 0);
    ------------------------ Receive Ports - RX AFE Ports ----------------------
    signal  gt0_gtprxn_i                    : std_logic;
    signal  gt0_gtprxp_i                    : std_logic;
    -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
    signal  gt0_rxcommadet_i                : std_logic;
    signal  gt0_rxmcommaalignen_i           : std_logic;
    signal  gt0_rxpcommaalignen_i           : std_logic;
    ------------ Receive Ports - RX Decision Feedback Equalizer(DFE) -----------
    signal  gt0_dmonitorout_i               : std_logic_vector(14 downto 0);
    -------------------- Receive Ports - RX Equailizer Ports -------------------
    signal  gt0_rxlpmhfhold_i               : std_logic;
    signal  gt0_rxlpmlfhold_i               : std_logic;
    --------------- Receive Ports - RX Fabric Output Control Ports -------------
    signal  gt0_rxoutclk_i                  : std_logic;
    signal  gt0_rxoutclkfabric_i            : std_logic;
    ------------- Receive Ports - RX Initialization and Reset Ports ------------
    signal  gt0_gtrxreset_i                 : std_logic;
    signal  gt0_rxlpmreset_i                : std_logic;
    -------------- Receive Ports -RX Initialization and Reset Ports ------------
    signal  gt0_rxresetdone_i               : std_logic;
    --------------------- TX Initialization and Reset Ports --------------------
    signal  gt0_gttxreset_i                 : std_logic;
    signal  gt0_txuserrdy_i                 : std_logic;
    ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
    signal  gt0_txdata_i                    : std_logic_vector(31 downto 0);
    ------------------ Transmit Ports - TX 8B/10B Encoder Ports ----------------
    signal  gt0_txcharisk_i                 : std_logic_vector(3 downto 0);
    --------------- Transmit Ports - TX Configurable Driver Ports --------------
    signal  gt0_gtptxn_i                    : std_logic;
    signal  gt0_gtptxp_i                    : std_logic;
    ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
    signal  gt0_txoutclk_i                  : std_logic;
    signal  gt0_txoutclkfabric_i            : std_logic;
    signal  gt0_txoutclkpcs_i               : std_logic;
    ------------- Transmit Ports - TX Initialization and Reset Ports -----------
    signal  gt0_txresetdone_i               : std_logic;

    --____________________________COMMON PORTS________________________________
   signal gt0_pll0reset_i  : std_logic;
   signal gt0_pll1reset_i  : std_logic;
   signal gt0_pll0reset_t  : std_logic;
   signal gt0_pll0pd_t  : std_logic;
   signal gt0_pll1pd_t  : std_logic;
   signal gt0_pll1reset_t  : std_logic;
         signal gt0_pll0outclk_i  : std_logic;
         signal gt0_pll0outrefclk_i  : std_logic;
         signal gt0_pll0lock_i  : std_logic;
         signal gt0_pll0refclklost_i  : std_logic;    
         signal gt0_pll1lock_i  : std_logic;
         signal gt0_pll1refclklost_i  : std_logic;    
         signal gt0_pll1outclk_i  : std_logic;
         signal gt0_pll1outrefclk_i  : std_logic;


    ------------------------------- Global Signals -----------------------------
    signal  gt0_tx_system_reset_c           : std_logic;
    signal  gt0_rx_system_reset_c           : std_logic;
    signal  tied_to_ground_i                : std_logic;
    signal  tied_to_ground_vec_i            : std_logic_vector(63 downto 0);
    signal  tied_to_vcc_i                   : std_logic;
    signal  tied_to_vcc_vec_i               : std_logic_vector(7 downto 0);
    signal  drpclk_in_i                     : std_logic;
    signal  sysclk_in_i                     : std_logic;
    signal  GTTXRESET_IN                    : std_logic;
    signal  GTRXRESET_IN                    : std_logic;
    signal  CPLLRESET_IN                    : std_logic;
    signal  QPLLRESET_IN                    : std_logic;

    attribute keep: string;
   ------------------------------- User Clocks ---------------------------------
    signal    gt0_txusrclk_i                  : std_logic; 
    signal    gt0_txusrclk2_i                 : std_logic; 
    signal    gt0_rxusrclk_i                  : std_logic; 
    signal    gt0_rxusrclk2_i                 : std_logic; 
    
    
    
    
    signal    gt0_txmmcm_lock_i               : std_logic;
    signal    gt0_txmmcm_reset_i              : std_logic;
    signal    gt0_rxmmcm_lock_i               : std_logic; 
    signal    gt0_rxmmcm_reset_i              : std_logic;
    ----------------------------- Reference Clocks ----------------------------
    
signal    q0_clk0_refclk_i                : std_logic;

signal commonreset_i : std_logic;

signal cpll_reset_pll0_q0_clk0_refclk_i : std_logic;
signal cpll_pd_pll0_q0_clk0_refclk_i : std_logic;


   attribute mark_debug                  : string;
   attribute mark_debug of SOFT_RESET_TX_IN : signal is "true";    
   attribute mark_debug of SOFT_RESET_RX_IN : signal is "true";
   attribute mark_debug of gt0_txmmcm_lock_i: signal is "true";
   attribute mark_debug of gt0_txmmcm_reset_i: signal is "true";
   attribute mark_debug of gt0_rxmmcm_lock_i: signal is "true";
   attribute mark_debug of gt0_rxmmcm_reset_i: signal is "true";
   attribute mark_debug of gt0_tx_fsm_reset_done_out: signal is "true";
   attribute mark_debug of gt0_rx_fsm_reset_done_out: signal is "true";
   attribute mark_debug of gt0_rxresetdone_out: signal is "true";
   attribute mark_debug of gt0_txresetdone_out: signal is "true";

   
   







--**************************** Main Body of Code *******************************
begin

refclk_out <= q0_clk0_refclk_i;

    --  Static signal Assigments
tied_to_ground_i                             <= '0';
tied_to_ground_vec_i                         <= x"0000000000000000";
tied_to_vcc_i                                <= '1';
tied_to_vcc_vec_i                            <= "11111111";

     GT0_TX_MMCM_LOCK_OUT <= gt0_txmmcm_lock_i;
    GT0_RX_MMCM_LOCK_OUT <= gt0_rxmmcm_lock_i;
 
    gt0_pll0reset_out <= commonreset_i or gt0_pll0reset_i;
     gt0_pll0outclk_out <= gt0_pll0outclk_i;
     gt0_pll0outrefclk_out <= gt0_pll0outrefclk_i;
     gt0_pll0reset_t <= commonreset_i or gt0_pll0reset_i or cpll_reset_pll0_q0_clk0_refclk_i;
     gt0_pll0pd_t <= cpll_pd_pll0_q0_clk0_refclk_i;
     gt0_pll0lock_out <= gt0_pll0lock_i;
     gt0_pll0refclklost_out <= gt0_pll0refclklost_i;    
     gt0_pll1outclk_out <= gt0_pll1outclk_i;
     gt0_pll1outrefclk_out <= gt0_pll1outrefclk_i;


 
      GT0_TXUSRCLK_OUT <= gt0_txusrclk_i; 
      GT0_TXUSRCLK2_OUT <= gt0_txusrclk2_i;
      GT0_RXUSRCLK_OUT <= gt0_rxusrclk_i;
      GT0_RXUSRCLK2_OUT <= gt0_rxusrclk2_i;


    
  
    gt_usrclk_source : kria_comm_GT_USRCLK_SOURCE
    port map
   (
 
        GT0_TXUSRCLK_OUT                =>      gt0_txusrclk_i,
        GT0_TXUSRCLK2_OUT               =>      gt0_txusrclk2_i,
        GT0_TXOUTCLK_IN                 =>      gt0_txoutclk_i,
        GT0_TXCLK_LOCK_OUT              =>      gt0_txmmcm_lock_i,
        GT0_TX_MMCM_RESET_IN            =>      gt0_txmmcm_reset_i,
        GT0_RXUSRCLK_OUT                =>      gt0_rxusrclk_i,
        GT0_RXUSRCLK2_OUT               =>      gt0_rxusrclk2_i,
        GT0_RXOUTCLK_IN                 =>      gt0_rxoutclk_i,
        GT0_RXCLK_LOCK_OUT              =>      gt0_rxmmcm_lock_i,
        GT0_RX_MMCM_RESET_IN            =>      gt0_rxmmcm_reset_i,
        Q0_CLK0_GTREFCLK_PAD_N_IN       =>      Q0_CLK0_GTREFCLK_PAD_N_IN,
        Q0_CLK0_GTREFCLK_PAD_P_IN       =>      Q0_CLK0_GTREFCLK_PAD_P_IN,
        Q0_CLK0_GTREFCLK_OUT            =>      q0_clk0_refclk_i

    );

sysclk_in_i <= sysclk_in;

  cpll_railing_pll0_q0_clk0_refclk_i : kria_comm_cpll_railing
  generic map(
           USE_BUFG       => 0
   ) 
   port map
   (
        cpll_reset_out => cpll_reset_pll0_q0_clk0_refclk_i,
        cpll_pd_out => cpll_pd_pll0_q0_clk0_refclk_i,
        refclk_out => open,
        refclk_in => q0_clk0_refclk_i 
); 



    common0_i:kria_comm_common 
  generic map
  (
   WRAPPER_SIM_GTRESET_SPEEDUP => EXAMPLE_SIM_GTRESET_SPEEDUP,
   SIM_PLL0REFCLK_SEL => "001",
   SIM_PLL1REFCLK_SEL => "001"
  )
 port map
   (
    PLL0OUTCLK_OUT => gt0_pll0outclk_i,
    PLL0OUTREFCLK_OUT => gt0_pll0outrefclk_i,
    PLL0LOCK_OUT => gt0_pll0lock_i,
    PLL0LOCKDETCLK_IN => sysclk_in_i,
    PLL0REFCLKLOST_OUT => gt0_pll0refclklost_i,    
    PLL0RESET_IN => gt0_pll0reset_t,
    PLL0REFCLKSEL_IN => "001",
    PLL0PD_IN => gt0_pll0pd_t,
    PLL1OUTCLK_OUT => gt0_pll1outclk_i,
    PLL1OUTREFCLK_OUT => gt0_pll1outrefclk_i,
    GTREFCLK0_IN => q0_clk0_refclk_i,

    GTREFCLK1_IN => tied_to_ground_i


);

    common_reset_i:kria_comm_common_reset 
   generic map 
   (
      STABLE_CLOCK_PERIOD =>STABLE_CLOCK_PERIOD        -- Period of the stable clock driving this state-machine, unit is [ns]
   )
   port map
   (    
      STABLE_CLOCK => sysclk_in_i,             --Stable Clock, either a stable clock from the PCB
      SOFT_RESET => soft_reset_tx_in,               --User Reset, can be pulled any time
      COMMON_RESET => commonreset_i              --Reset QPLL
   );


    kria_comm_init_i : kria_comm
    port map
    (
        sysclk_in                       =>      sysclk_in_i,
        soft_reset_tx_in                =>      SOFT_RESET_TX_IN,
        soft_reset_rx_in                =>      SOFT_RESET_RX_IN,
        dont_reset_on_data_error_in     =>      DONT_RESET_ON_DATA_ERROR_IN,
        gt0_tx_mmcm_lock_in             =>      gt0_txmmcm_lock_i,
        gt0_tx_mmcm_reset_out           =>      gt0_txmmcm_reset_i,
        gt0_rx_mmcm_lock_in             =>      gt0_rxmmcm_lock_i,
        gt0_rx_mmcm_reset_out           =>      gt0_rxmmcm_reset_i,
        gt0_drp_busy_out                =>      open,
        gt0_tx_fsm_reset_done_out       =>      gt0_tx_fsm_reset_done_out,
        gt0_rx_fsm_reset_done_out       =>      gt0_rx_fsm_reset_done_out,
        gt0_data_valid_in               =>      gt0_data_valid_in,

        --_____________________________________________________________________
        --_____________________________________________________________________
        --GT0  (X0Y0)

        ---------------------------- Channel - DRP Ports  --------------------------
        gt0_drpaddr_in                  =>      gt0_drpaddr_in,
        gt0_drpclk_in                   =>      sysclk_in_i,
        gt0_drpdi_in                    =>      gt0_drpdi_in,
        gt0_drpdo_out                   =>      gt0_drpdo_out,
        gt0_drpen_in                    =>      gt0_drpen_in,
        gt0_drprdy_out                  =>      gt0_drprdy_out,
        gt0_drpwe_in                    =>      gt0_drpwe_in,
        --------------------- RX Initialization and Reset Ports --------------------
        gt0_eyescanreset_in             =>      gt0_eyescanreset_in,
        gt0_rxuserrdy_in                =>      gt0_rxuserrdy_in,
        -------------------------- RX Margin Analysis Ports ------------------------
        gt0_eyescandataerror_out        =>      gt0_eyescandataerror_out,
        gt0_eyescantrigger_in           =>      gt0_eyescantrigger_in,
        ------------------ Receive Ports - FPGA RX Interface Ports -----------------
        gt0_rxdata_out                  =>      gt0_rxdata_out,
        gt0_rxusrclk_in                 =>      gt0_rxusrclk_i,
        gt0_rxusrclk2_in                =>      gt0_rxusrclk2_i,
        ------------------ Receive Ports - RX 8B/10B Decoder Ports -----------------
        gt0_rxchariscomma_out           =>      gt0_rxchariscomma_out,
        gt0_rxcharisk_out               =>      gt0_rxcharisk_out,
        gt0_rxdisperr_out               =>      gt0_rxdisperr_out,
        gt0_rxnotintable_out            =>      gt0_rxnotintable_out,
        ------------------------ Receive Ports - RX AFE Ports ----------------------
        gt0_gtprxn_in                   =>      gt0_gtprxn_in,
        gt0_gtprxp_in                   =>      gt0_gtprxp_in,
        -------------- Receive Ports - RX Byte and Word Alignment Ports ------------
        gt0_rxcommadet_out              =>      gt0_rxcommadet_out,
        gt0_rxmcommaalignen_in          =>      gt0_rxmcommaalignen_in,
        gt0_rxpcommaalignen_in          =>      gt0_rxpcommaalignen_in,
        ------------ Receive Ports - RX Decision Feedback Equalizer(DFE) -----------
        gt0_dmonitorout_out             =>      gt0_dmonitorout_out,
        -------------------- Receive Ports - RX Equailizer Ports -------------------
        gt0_rxlpmhfhold_in              =>      gt0_rxlpmhfhold_in,
        gt0_rxlpmlfhold_in              =>      gt0_rxlpmlfhold_in,
        --------------- Receive Ports - RX Fabric Output Control Ports -------------
        gt0_rxoutclk_out                =>      gt0_rxoutclk_i,
        gt0_rxoutclkfabric_out          =>      gt0_rxoutclkfabric_out,
        ------------- Receive Ports - RX Initialization and Reset Ports ------------
        gt0_gtrxreset_in                =>      gt0_gtrxreset_in,
        gt0_rxlpmreset_in               =>      gt0_rxlpmreset_in,
        ----------------- Receive Ports - RX Polarity Control Ports ----------------
        gt0_rxpolarity_in               =>      '1',         
            
        -------------- Receive Ports -RX Initialization and Reset Ports ------------
        gt0_rxresetdone_out             =>      gt0_rxresetdone_out,
        --------------------- TX Initialization and Reset Ports --------------------
        gt0_gttxreset_in                =>      gt0_gttxreset_in,
        gt0_txuserrdy_in                =>      gt0_txuserrdy_in,
        ------------------ Transmit Ports - FPGA TX Interface Ports ----------------
        gt0_txdata_in                   =>      gt0_txdata_in,
        gt0_txusrclk_in                 =>      gt0_txusrclk_i,
        gt0_txusrclk2_in                =>      gt0_txusrclk2_i,
        ------------------ Transmit Ports - TX 8B/10B Encoder Ports ----------------
        gt0_txcharisk_in                =>      gt0_txcharisk_in,
        --------------- Transmit Ports - TX Configurable Driver Ports --------------
        gt0_gtptxn_out                  =>      gt0_gtptxn_out,
        gt0_gtptxp_out                  =>      gt0_gtptxp_out,
        ----------- Transmit Ports - TX Fabric Clock Output Control Ports ----------
        gt0_txoutclk_out                =>      gt0_txoutclk_i,
        gt0_txoutclkfabric_out          =>      gt0_txoutclkfabric_out,
        gt0_txoutclkpcs_out             =>      gt0_txoutclkpcs_out,
        ------------- Transmit Ports - TX Initialization and Reset Ports -----------
        gt0_txresetdone_out             =>      gt0_txresetdone_out,

        gt0_pll0outclk_in               =>      gt0_pll0outclk_i,
        gt0_pll0outrefclk_in            =>      gt0_pll0outrefclk_i,
        gt0_pll0reset_out               =>      gt0_pll0reset_i,
        gt0_pll0lock_in                 =>      gt0_pll0lock_i,
        gt0_pll0refclklost_in           =>      gt0_pll0refclklost_i,    
        gt0_pll1outclk_in               =>      gt0_pll1outclk_i,
        gt0_pll1outrefclk_in            =>      gt0_pll1outrefclk_i
    );



end RTL;
